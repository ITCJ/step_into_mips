`include "defines.v"

module mem(
    input rst,

    input rw_i,
    input wreg_i,
    input wdata_i,

    output reg rw_o,
    output reg wreg_o,
    output reg wdata_o
);

endmodule