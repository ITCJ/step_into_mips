`include "defines.v"

module regfile(
    input 
);