module pc_reg(
    input rst,
    input clk,

    output reg pc,
    output reg ce
    );


endmodule
